-- Bibliotecas
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

--Entidad

entity Entidad_6 is

--Declaracion de puertos

port(
	--Entradas A,B y C
	Entradas: in std_LOGIC_1164
	
)